module display(
    input logic [11 : 0] sum_result,
    output logic [6 : 0] units,
    output logic [6 : 0] tens,
    output logic [6 : 0] hundreds,
    output logic [6 : 0] thousands
);

    //Almacena temporalmente cada dígito
    logic [3:0] units_digit;
    logic [3:0] tens_digit;
    logic [3:0] hundreds_digit;
    logic [3:0] thousands_digit;





endmodule